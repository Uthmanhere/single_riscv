module our;
	initial begin $display("Hello world"); $finish; end
endmodule

