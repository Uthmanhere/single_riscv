module alu_cu (
	input	[2:0]	funct3,
	input			funct7,
	input	[1:0]	aluOp_cu
)

	always_comb begin
		case (aluOp_cu)
			00 :
			01 :
			10 :
			11 :

	end

endmodule
