module alu (

		input [31:0]	r1,
		input [31:0]	r2,
		input [2:0]		alu_ctrl,
		output			zero,
		output [31:0]	aluOut

	);

	


endmodule
