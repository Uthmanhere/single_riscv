`include "alu.sv"
`include "pc.sv"
`include "dataMem.sv"
`include "instMem.sv"
`include "regfile.sv"

module rv32i (

	input	clk

)

	


endmodule
