module alu_cu (
	input	[2:0]	funct3,
	input			funct7,
	input	[1:0]	aluOp_cu
)



endmodule
